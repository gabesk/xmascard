`timescale 1ns / 1ps

//
// Validates that updating a pattern works according to design.
//


// In testing on the hardware, PuTTY was having trouble reliably sending and
// receiving the lowercase letter 'a'. Nothing else; the test data here worked
// fine. So this variation attempts to figure out why.
// Wait a random amount of time, then send 'a', repeatedly over and over. If the
// receiver ever receives something other than 'a' back, assert.

module test;

    // Inputs
    reg clk = 0;
    reg rx = 1; // RS-232 idle condition is logic high
    reg xmit = 0;
    reg recv = 0;
    reg write_complete_received = 0;
    reg test_step_complete = 0;

    integer i = 0;
    integer j = 0;
    integer random_delay;
    reg [7:0] received_byte = 0;

    reg [7:0] test_send_vector [0:576];
    integer test_send_vector_len = 576;
    reg [7:0] test_receive_vector [0:384];
    integer test_receive_vector_len = 384;
    
    initial begin
        test_send_vector[0]  = "i";
        test_send_vector[1]  = 8'h0;
        test_send_vector[2]  = 8'h0;
        test_send_vector[3]  = "i";
        test_send_vector[4]  = 8'h0;
        test_send_vector[5]  = 8'h1;
        test_send_vector[6]  = "i";
        test_send_vector[7]  = 8'h0;
        test_send_vector[8]  = 8'h2;
        test_send_vector[9]  = "i";
        test_send_vector[10]  = 8'h0;
        test_send_vector[11]  = 8'h3;
        test_send_vector[12]  = "i";
        test_send_vector[13]  = 8'h0;
        test_send_vector[14]  = 8'h4;
        test_send_vector[15]  = "i";
        test_send_vector[16]  = 8'h0;
        test_send_vector[17]  = 8'h5;
        test_send_vector[18]  = "i";
        test_send_vector[19]  = 8'h0;
        test_send_vector[20]  = 8'h6;
        test_send_vector[21]  = "i";
        test_send_vector[22]  = 8'h0;
        test_send_vector[23]  = 8'h7;
        test_send_vector[24]  = "i";
        test_send_vector[25]  = 8'h1;
        test_send_vector[26]  = 8'h0;
        test_send_vector[27]  = "i";
        test_send_vector[28]  = 8'h1;
        test_send_vector[29]  = 8'h1;
        test_send_vector[30]  = "i";
        test_send_vector[31]  = 8'h1;
        test_send_vector[32]  = 8'h2;
        test_send_vector[33]  = "i";
        test_send_vector[34]  = 8'h1;
        test_send_vector[35]  = 8'h3;
        test_send_vector[36]  = "i";
        test_send_vector[37]  = 8'h1;
        test_send_vector[38]  = 8'h4;
        test_send_vector[39]  = "i";
        test_send_vector[40]  = 8'h1;
        test_send_vector[41]  = 8'h5;
        test_send_vector[42]  = "i";
        test_send_vector[43]  = 8'h1;
        test_send_vector[44]  = 8'h6;
        test_send_vector[45]  = "i";
        test_send_vector[46]  = 8'h1;
        test_send_vector[47]  = 8'h7;
        test_send_vector[48]  = "i";
        test_send_vector[49]  = 8'h2;
        test_send_vector[50]  = 8'h0;
        test_send_vector[51]  = "i";
        test_send_vector[52]  = 8'h2;
        test_send_vector[53]  = 8'h1;
        test_send_vector[54]  = "i";
        test_send_vector[55]  = 8'h2;
        test_send_vector[56]  = 8'h2;
        test_send_vector[57]  = "i";
        test_send_vector[58]  = 8'h2;
        test_send_vector[59]  = 8'h3;
        test_send_vector[60]  = "i";
        test_send_vector[61]  = 8'h2;
        test_send_vector[62]  = 8'h4;
        test_send_vector[63]  = "i";
        test_send_vector[64]  = 8'h2;
        test_send_vector[65]  = 8'h5;
        test_send_vector[66]  = "i";
        test_send_vector[67]  = 8'h2;
        test_send_vector[68]  = 8'h6;
        test_send_vector[69]  = "i";
        test_send_vector[70]  = 8'h2;
        test_send_vector[71]  = 8'h7;
        test_send_vector[72]  = "i";
        test_send_vector[73]  = 8'h3;
        test_send_vector[74]  = 8'h0;
        test_send_vector[75]  = "i";
        test_send_vector[76]  = 8'h3;
        test_send_vector[77]  = 8'h1;
        test_send_vector[78]  = "i";
        test_send_vector[79]  = 8'h3;
        test_send_vector[80]  = 8'h2;
        test_send_vector[81]  = "i";
        test_send_vector[82]  = 8'h3;
        test_send_vector[83]  = 8'h3;
        test_send_vector[84]  = "i";
        test_send_vector[85]  = 8'h3;
        test_send_vector[86]  = 8'h4;
        test_send_vector[87]  = "i";
        test_send_vector[88]  = 8'h3;
        test_send_vector[89]  = 8'h5;
        test_send_vector[90]  = "i";
        test_send_vector[91]  = 8'h3;
        test_send_vector[92]  = 8'h6;
        test_send_vector[93]  = "i";
        test_send_vector[94]  = 8'h3;
        test_send_vector[95]  = 8'h7;
        test_send_vector[96]  = "i";
        test_send_vector[97]  = 8'h4;
        test_send_vector[98]  = 8'h0;
        test_send_vector[99]  = "i";
        test_send_vector[100]  = 8'h4;
        test_send_vector[101]  = 8'h1;
        test_send_vector[102]  = "i";
        test_send_vector[103]  = 8'h4;
        test_send_vector[104]  = 8'h2;
        test_send_vector[105]  = "i";
        test_send_vector[106]  = 8'h4;
        test_send_vector[107]  = 8'h3;
        test_send_vector[108]  = "i";
        test_send_vector[109]  = 8'h4;
        test_send_vector[110]  = 8'h4;
        test_send_vector[111]  = "i";
        test_send_vector[112]  = 8'h4;
        test_send_vector[113]  = 8'h5;
        test_send_vector[114]  = "i";
        test_send_vector[115]  = 8'h4;
        test_send_vector[116]  = 8'h6;
        test_send_vector[117]  = "i";
        test_send_vector[118]  = 8'h4;
        test_send_vector[119]  = 8'h7;
        test_send_vector[120]  = "i";
        test_send_vector[121]  = 8'h5;
        test_send_vector[122]  = 8'h0;
        test_send_vector[123]  = "i";
        test_send_vector[124]  = 8'h5;
        test_send_vector[125]  = 8'h1;
        test_send_vector[126]  = "i";
        test_send_vector[127]  = 8'h5;
        test_send_vector[128]  = 8'h2;
        test_send_vector[129]  = "i";
        test_send_vector[130]  = 8'h5;
        test_send_vector[131]  = 8'h3;
        test_send_vector[132]  = "i";
        test_send_vector[133]  = 8'h5;
        test_send_vector[134]  = 8'h4;
        test_send_vector[135]  = "i";
        test_send_vector[136]  = 8'h5;
        test_send_vector[137]  = 8'h5;
        test_send_vector[138]  = "i";
        test_send_vector[139]  = 8'h5;
        test_send_vector[140]  = 8'h6;
        test_send_vector[141]  = "i";
        test_send_vector[142]  = 8'h5;
        test_send_vector[143]  = 8'h7;
        test_send_vector[144]  = "i";
        test_send_vector[145]  = 8'h6;
        test_send_vector[146]  = 8'h0;
        test_send_vector[147]  = "i";
        test_send_vector[148]  = 8'h6;
        test_send_vector[149]  = 8'h1;
        test_send_vector[150]  = "i";
        test_send_vector[151]  = 8'h6;
        test_send_vector[152]  = 8'h2;
        test_send_vector[153]  = "i";
        test_send_vector[154]  = 8'h6;
        test_send_vector[155]  = 8'h3;
        test_send_vector[156]  = "i";
        test_send_vector[157]  = 8'h6;
        test_send_vector[158]  = 8'h4;
        test_send_vector[159]  = "i";
        test_send_vector[160]  = 8'h6;
        test_send_vector[161]  = 8'h5;
        test_send_vector[162]  = "i";
        test_send_vector[163]  = 8'h6;
        test_send_vector[164]  = 8'h6;
        test_send_vector[165]  = "i";
        test_send_vector[166]  = 8'h6;
        test_send_vector[167]  = 8'h7;
        test_send_vector[168]  = "i";
        test_send_vector[169]  = 8'h7;
        test_send_vector[170]  = 8'h0;
        test_send_vector[171]  = "i";
        test_send_vector[172]  = 8'h7;
        test_send_vector[173]  = 8'h1;
        test_send_vector[174]  = "i";
        test_send_vector[175]  = 8'h7;
        test_send_vector[176]  = 8'h2;
        test_send_vector[177]  = "i";
        test_send_vector[178]  = 8'h7;
        test_send_vector[179]  = 8'h3;
        test_send_vector[180]  = "i";
        test_send_vector[181]  = 8'h7;
        test_send_vector[182]  = 8'h4;
        test_send_vector[183]  = "i";
        test_send_vector[184]  = 8'h7;
        test_send_vector[185]  = 8'h5;
        test_send_vector[186]  = "i";
        test_send_vector[187]  = 8'h7;
        test_send_vector[188]  = 8'h6;
        test_send_vector[189]  = "i";
        test_send_vector[190]  = 8'h7;
        test_send_vector[191]  = 8'h7;
        test_send_vector[192]  = "i";
        test_send_vector[193]  = 8'h8;
        test_send_vector[194]  = 8'h0;
        test_send_vector[195]  = "i";
        test_send_vector[196]  = 8'h8;
        test_send_vector[197]  = 8'h1;
        test_send_vector[198]  = "i";
        test_send_vector[199]  = 8'h8;
        test_send_vector[200]  = 8'h2;
        test_send_vector[201]  = "i";
        test_send_vector[202]  = 8'h8;
        test_send_vector[203]  = 8'h3;
        test_send_vector[204]  = "i";
        test_send_vector[205]  = 8'h8;
        test_send_vector[206]  = 8'h4;
        test_send_vector[207]  = "i";
        test_send_vector[208]  = 8'h8;
        test_send_vector[209]  = 8'h5;
        test_send_vector[210]  = "i";
        test_send_vector[211]  = 8'h8;
        test_send_vector[212]  = 8'h6;
        test_send_vector[213]  = "i";
        test_send_vector[214]  = 8'h8;
        test_send_vector[215]  = 8'h7;
        test_send_vector[216]  = "i";
        test_send_vector[217]  = 8'h9;
        test_send_vector[218]  = 8'h0;
        test_send_vector[219]  = "i";
        test_send_vector[220]  = 8'h9;
        test_send_vector[221]  = 8'h1;
        test_send_vector[222]  = "i";
        test_send_vector[223]  = 8'h9;
        test_send_vector[224]  = 8'h2;
        test_send_vector[225]  = "i";
        test_send_vector[226]  = 8'h9;
        test_send_vector[227]  = 8'h3;
        test_send_vector[228]  = "i";
        test_send_vector[229]  = 8'h9;
        test_send_vector[230]  = 8'h4;
        test_send_vector[231]  = "i";
        test_send_vector[232]  = 8'h9;
        test_send_vector[233]  = 8'h5;
        test_send_vector[234]  = "i";
        test_send_vector[235]  = 8'h9;
        test_send_vector[236]  = 8'h6;
        test_send_vector[237]  = "i";
        test_send_vector[238]  = 8'h9;
        test_send_vector[239]  = 8'h7;
        test_send_vector[240]  = "i";
        test_send_vector[241]  = 8'ha;
        test_send_vector[242]  = 8'h0;
        test_send_vector[243]  = "i";
        test_send_vector[244]  = 8'ha;
        test_send_vector[245]  = 8'h1;
        test_send_vector[246]  = "i";
        test_send_vector[247]  = 8'ha;
        test_send_vector[248]  = 8'h2;
        test_send_vector[249]  = "i";
        test_send_vector[250]  = 8'ha;
        test_send_vector[251]  = 8'h3;
        test_send_vector[252]  = "i";
        test_send_vector[253]  = 8'ha;
        test_send_vector[254]  = 8'h4;
        test_send_vector[255]  = "i";
        test_send_vector[256]  = 8'ha;
        test_send_vector[257]  = 8'h5;
        test_send_vector[258]  = "i";
        test_send_vector[259]  = 8'ha;
        test_send_vector[260]  = 8'h6;
        test_send_vector[261]  = "i";
        test_send_vector[262]  = 8'ha;
        test_send_vector[263]  = 8'h7;
        test_send_vector[264]  = "i";
        test_send_vector[265]  = 8'hb;
        test_send_vector[266]  = 8'h0;
        test_send_vector[267]  = "i";
        test_send_vector[268]  = 8'hb;
        test_send_vector[269]  = 8'h1;
        test_send_vector[270]  = "i";
        test_send_vector[271]  = 8'hb;
        test_send_vector[272]  = 8'h2;
        test_send_vector[273]  = "i";
        test_send_vector[274]  = 8'hb;
        test_send_vector[275]  = 8'h3;
        test_send_vector[276]  = "i";
        test_send_vector[277]  = 8'hb;
        test_send_vector[278]  = 8'h4;
        test_send_vector[279]  = "i";
        test_send_vector[280]  = 8'hb;
        test_send_vector[281]  = 8'h5;
        test_send_vector[282]  = "i";
        test_send_vector[283]  = 8'hb;
        test_send_vector[284]  = 8'h6;
        test_send_vector[285]  = "i";
        test_send_vector[286]  = 8'hb;
        test_send_vector[287]  = 8'h7;
        test_send_vector[288]  = "i";
        test_send_vector[289]  = 8'hc;
        test_send_vector[290]  = 8'h0;
        test_send_vector[291]  = "i";
        test_send_vector[292]  = 8'hc;
        test_send_vector[293]  = 8'h1;
        test_send_vector[294]  = "i";
        test_send_vector[295]  = 8'hc;
        test_send_vector[296]  = 8'h2;
        test_send_vector[297]  = "i";
        test_send_vector[298]  = 8'hc;
        test_send_vector[299]  = 8'h3;
        test_send_vector[300]  = "i";
        test_send_vector[301]  = 8'hc;
        test_send_vector[302]  = 8'h4;
        test_send_vector[303]  = "i";
        test_send_vector[304]  = 8'hc;
        test_send_vector[305]  = 8'h5;
        test_send_vector[306]  = "i";
        test_send_vector[307]  = 8'hc;
        test_send_vector[308]  = 8'h6;
        test_send_vector[309]  = "i";
        test_send_vector[310]  = 8'hc;
        test_send_vector[311]  = 8'h7;
        test_send_vector[312]  = "i";
        test_send_vector[313]  = 8'hd;
        test_send_vector[314]  = 8'h0;
        test_send_vector[315]  = "i";
        test_send_vector[316]  = 8'hd;
        test_send_vector[317]  = 8'h1;
        test_send_vector[318]  = "i";
        test_send_vector[319]  = 8'hd;
        test_send_vector[320]  = 8'h2;
        test_send_vector[321]  = "i";
        test_send_vector[322]  = 8'hd;
        test_send_vector[323]  = 8'h3;
        test_send_vector[324]  = "i";
        test_send_vector[325]  = 8'hd;
        test_send_vector[326]  = 8'h4;
        test_send_vector[327]  = "i";
        test_send_vector[328]  = 8'hd;
        test_send_vector[329]  = 8'h5;
        test_send_vector[330]  = "i";
        test_send_vector[331]  = 8'hd;
        test_send_vector[332]  = 8'h6;
        test_send_vector[333]  = "i";
        test_send_vector[334]  = 8'hd;
        test_send_vector[335]  = 8'h7;
        test_send_vector[336]  = "i";
        test_send_vector[337]  = 8'he;
        test_send_vector[338]  = 8'h0;
        test_send_vector[339]  = "i";
        test_send_vector[340]  = 8'he;
        test_send_vector[341]  = 8'h1;
        test_send_vector[342]  = "i";
        test_send_vector[343]  = 8'he;
        test_send_vector[344]  = 8'h2;
        test_send_vector[345]  = "i";
        test_send_vector[346]  = 8'he;
        test_send_vector[347]  = 8'h3;
        test_send_vector[348]  = "i";
        test_send_vector[349]  = 8'he;
        test_send_vector[350]  = 8'h4;
        test_send_vector[351]  = "i";
        test_send_vector[352]  = 8'he;
        test_send_vector[353]  = 8'h5;
        test_send_vector[354]  = "i";
        test_send_vector[355]  = 8'he;
        test_send_vector[356]  = 8'h6;
        test_send_vector[357]  = "i";
        test_send_vector[358]  = 8'he;
        test_send_vector[359]  = 8'h7;
        test_send_vector[360]  = "i";
        test_send_vector[361]  = 8'hf;
        test_send_vector[362]  = 8'h0;
        test_send_vector[363]  = "i";
        test_send_vector[364]  = 8'hf;
        test_send_vector[365]  = 8'h1;
        test_send_vector[366]  = "i";
        test_send_vector[367]  = 8'hf;
        test_send_vector[368]  = 8'h2;
        test_send_vector[369]  = "i";
        test_send_vector[370]  = 8'hf;
        test_send_vector[371]  = 8'h3;
        test_send_vector[372]  = "i";
        test_send_vector[373]  = 8'hf;
        test_send_vector[374]  = 8'h4;
        test_send_vector[375]  = "i";
        test_send_vector[376]  = 8'hf;
        test_send_vector[377]  = 8'h5;
        test_send_vector[378]  = "i";
        test_send_vector[379]  = 8'hf;
        test_send_vector[380]  = 8'h6;
        test_send_vector[381]  = "i";
        test_send_vector[382]  = 8'hf;
        test_send_vector[383]  = 8'h7;
        test_send_vector[384]  = "i";
        test_send_vector[385]  = 8'h10;
        test_send_vector[386]  = 8'h0;
        test_send_vector[387]  = "i";
        test_send_vector[388]  = 8'h10;
        test_send_vector[389]  = 8'h1;
        test_send_vector[390]  = "i";
        test_send_vector[391]  = 8'h10;
        test_send_vector[392]  = 8'h2;
        test_send_vector[393]  = "i";
        test_send_vector[394]  = 8'h10;
        test_send_vector[395]  = 8'h3;
        test_send_vector[396]  = "i";
        test_send_vector[397]  = 8'h10;
        test_send_vector[398]  = 8'h4;
        test_send_vector[399]  = "i";
        test_send_vector[400]  = 8'h10;
        test_send_vector[401]  = 8'h5;
        test_send_vector[402]  = "i";
        test_send_vector[403]  = 8'h10;
        test_send_vector[404]  = 8'h6;
        test_send_vector[405]  = "i";
        test_send_vector[406]  = 8'h10;
        test_send_vector[407]  = 8'h7;
        test_send_vector[408]  = "i";
        test_send_vector[409]  = 8'h11;
        test_send_vector[410]  = 8'h0;
        test_send_vector[411]  = "i";
        test_send_vector[412]  = 8'h11;
        test_send_vector[413]  = 8'h1;
        test_send_vector[414]  = "i";
        test_send_vector[415]  = 8'h11;
        test_send_vector[416]  = 8'h2;
        test_send_vector[417]  = "i";
        test_send_vector[418]  = 8'h11;
        test_send_vector[419]  = 8'h3;
        test_send_vector[420]  = "i";
        test_send_vector[421]  = 8'h11;
        test_send_vector[422]  = 8'h4;
        test_send_vector[423]  = "i";
        test_send_vector[424]  = 8'h11;
        test_send_vector[425]  = 8'h5;
        test_send_vector[426]  = "i";
        test_send_vector[427]  = 8'h11;
        test_send_vector[428]  = 8'h6;
        test_send_vector[429]  = "i";
        test_send_vector[430]  = 8'h11;
        test_send_vector[431]  = 8'h7;
        test_send_vector[432]  = "i";
        test_send_vector[433]  = 8'h12;
        test_send_vector[434]  = 8'h0;
        test_send_vector[435]  = "i";
        test_send_vector[436]  = 8'h12;
        test_send_vector[437]  = 8'h1;
        test_send_vector[438]  = "i";
        test_send_vector[439]  = 8'h12;
        test_send_vector[440]  = 8'h2;
        test_send_vector[441]  = "i";
        test_send_vector[442]  = 8'h12;
        test_send_vector[443]  = 8'h3;
        test_send_vector[444]  = "i";
        test_send_vector[445]  = 8'h12;
        test_send_vector[446]  = 8'h4;
        test_send_vector[447]  = "i";
        test_send_vector[448]  = 8'h12;
        test_send_vector[449]  = 8'h5;
        test_send_vector[450]  = "i";
        test_send_vector[451]  = 8'h12;
        test_send_vector[452]  = 8'h6;
        test_send_vector[453]  = "i";
        test_send_vector[454]  = 8'h12;
        test_send_vector[455]  = 8'h7;
        test_send_vector[456]  = "i";
        test_send_vector[457]  = 8'h13;
        test_send_vector[458]  = 8'h0;
        test_send_vector[459]  = "i";
        test_send_vector[460]  = 8'h13;
        test_send_vector[461]  = 8'h1;
        test_send_vector[462]  = "i";
        test_send_vector[463]  = 8'h13;
        test_send_vector[464]  = 8'h2;
        test_send_vector[465]  = "i";
        test_send_vector[466]  = 8'h13;
        test_send_vector[467]  = 8'h3;
        test_send_vector[468]  = "i";
        test_send_vector[469]  = 8'h13;
        test_send_vector[470]  = 8'h4;
        test_send_vector[471]  = "i";
        test_send_vector[472]  = 8'h13;
        test_send_vector[473]  = 8'h5;
        test_send_vector[474]  = "i";
        test_send_vector[475]  = 8'h13;
        test_send_vector[476]  = 8'h6;
        test_send_vector[477]  = "i";
        test_send_vector[478]  = 8'h13;
        test_send_vector[479]  = 8'h7;
        test_send_vector[480]  = "i";
        test_send_vector[481]  = 8'h14;
        test_send_vector[482]  = 8'h0;
        test_send_vector[483]  = "i";
        test_send_vector[484]  = 8'h14;
        test_send_vector[485]  = 8'h1;
        test_send_vector[486]  = "i";
        test_send_vector[487]  = 8'h14;
        test_send_vector[488]  = 8'h2;
        test_send_vector[489]  = "i";
        test_send_vector[490]  = 8'h14;
        test_send_vector[491]  = 8'h3;
        test_send_vector[492]  = "i";
        test_send_vector[493]  = 8'h14;
        test_send_vector[494]  = 8'h4;
        test_send_vector[495]  = "i";
        test_send_vector[496]  = 8'h14;
        test_send_vector[497]  = 8'h5;
        test_send_vector[498]  = "i";
        test_send_vector[499]  = 8'h14;
        test_send_vector[500]  = 8'h6;
        test_send_vector[501]  = "i";
        test_send_vector[502]  = 8'h14;
        test_send_vector[503]  = 8'h7;
        test_send_vector[504]  = "i";
        test_send_vector[505]  = 8'h15;
        test_send_vector[506]  = 8'h0;
        test_send_vector[507]  = "i";
        test_send_vector[508]  = 8'h15;
        test_send_vector[509]  = 8'h1;
        test_send_vector[510]  = "i";
        test_send_vector[511]  = 8'h15;
        test_send_vector[512]  = 8'h2;
        test_send_vector[513]  = "i";
        test_send_vector[514]  = 8'h15;
        test_send_vector[515]  = 8'h3;
        test_send_vector[516]  = "i";
        test_send_vector[517]  = 8'h15;
        test_send_vector[518]  = 8'h4;
        test_send_vector[519]  = "i";
        test_send_vector[520]  = 8'h15;
        test_send_vector[521]  = 8'h5;
        test_send_vector[522]  = "i";
        test_send_vector[523]  = 8'h15;
        test_send_vector[524]  = 8'h6;
        test_send_vector[525]  = "i";
        test_send_vector[526]  = 8'h15;
        test_send_vector[527]  = 8'h7;
        test_send_vector[528]  = "i";
        test_send_vector[529]  = 8'h16;
        test_send_vector[530]  = 8'h0;
        test_send_vector[531]  = "i";
        test_send_vector[532]  = 8'h16;
        test_send_vector[533]  = 8'h1;
        test_send_vector[534]  = "i";
        test_send_vector[535]  = 8'h16;
        test_send_vector[536]  = 8'h2;
        test_send_vector[537]  = "i";
        test_send_vector[538]  = 8'h16;
        test_send_vector[539]  = 8'h3;
        test_send_vector[540]  = "i";
        test_send_vector[541]  = 8'h16;
        test_send_vector[542]  = 8'h4;
        test_send_vector[543]  = "i";
        test_send_vector[544]  = 8'h16;
        test_send_vector[545]  = 8'h5;
        test_send_vector[546]  = "i";
        test_send_vector[547]  = 8'h16;
        test_send_vector[548]  = 8'h6;
        test_send_vector[549]  = "i";
        test_send_vector[550]  = 8'h16;
        test_send_vector[551]  = 8'h7;
        test_send_vector[552]  = "i";
        test_send_vector[553]  = 8'h17;
        test_send_vector[554]  = 8'h0;
        test_send_vector[555]  = "i";
        test_send_vector[556]  = 8'h17;
        test_send_vector[557]  = 8'h1;
        test_send_vector[558]  = "i";
        test_send_vector[559]  = 8'h17;
        test_send_vector[560]  = 8'h2;
        test_send_vector[561]  = "i";
        test_send_vector[562]  = 8'h17;
        test_send_vector[563]  = 8'h3;
        test_send_vector[564]  = "i";
        test_send_vector[565]  = 8'h17;
        test_send_vector[566]  = 8'h4;
        test_send_vector[567]  = "i";
        test_send_vector[568]  = 8'h17;
        test_send_vector[569]  = 8'h5;
        test_send_vector[570]  = "i";
        test_send_vector[571]  = 8'h17;
        test_send_vector[572]  = 8'h6;
        test_send_vector[573]  = "i";
        test_send_vector[574]  = 8'h17;
        test_send_vector[575]  = 8'h7;
        test_receive_vector[0]  = 8'h0;
        test_receive_vector[1]  = 8'h0;
        test_receive_vector[2]  = 8'h0;
        test_receive_vector[3]  = 8'h1;
        test_receive_vector[4]  = 8'h0;
        test_receive_vector[5]  = 8'h2;
        test_receive_vector[6]  = 8'h0;
        test_receive_vector[7]  = 8'h3;
        test_receive_vector[8]  = 8'h0;
        test_receive_vector[9]  = 8'h4;
        test_receive_vector[10]  = 8'h0;
        test_receive_vector[11]  = 8'h5;
        test_receive_vector[12]  = 8'h0;
        test_receive_vector[13]  = 8'h6;
        test_receive_vector[14]  = 8'h0;
        test_receive_vector[15]  = 8'h7;
        test_receive_vector[16]  = 8'h1;
        test_receive_vector[17]  = 8'h0;
        test_receive_vector[18]  = 8'h1;
        test_receive_vector[19]  = 8'h1;
        test_receive_vector[20]  = 8'h1;
        test_receive_vector[21]  = 8'h2;
        test_receive_vector[22]  = 8'h1;
        test_receive_vector[23]  = 8'h3;
        test_receive_vector[24]  = 8'h1;
        test_receive_vector[25]  = 8'h4;
        test_receive_vector[26]  = 8'h1;
        test_receive_vector[27]  = 8'h5;
        test_receive_vector[28]  = 8'h1;
        test_receive_vector[29]  = 8'h6;
        test_receive_vector[30]  = 8'h1;
        test_receive_vector[31]  = 8'h7;
        test_receive_vector[32]  = 8'h2;
        test_receive_vector[33]  = 8'h0;
        test_receive_vector[34]  = 8'h2;
        test_receive_vector[35]  = 8'h1;
        test_receive_vector[36]  = 8'h2;
        test_receive_vector[37]  = 8'h2;
        test_receive_vector[38]  = 8'h2;
        test_receive_vector[39]  = 8'h3;
        test_receive_vector[40]  = 8'h2;
        test_receive_vector[41]  = 8'h4;
        test_receive_vector[42]  = 8'h2;
        test_receive_vector[43]  = 8'h5;
        test_receive_vector[44]  = 8'h2;
        test_receive_vector[45]  = 8'h6;
        test_receive_vector[46]  = 8'h2;
        test_receive_vector[47]  = 8'h7;
        test_receive_vector[48]  = 8'h3;
        test_receive_vector[49]  = 8'h0;
        test_receive_vector[50]  = 8'h3;
        test_receive_vector[51]  = 8'h1;
        test_receive_vector[52]  = 8'h3;
        test_receive_vector[53]  = 8'h2;
        test_receive_vector[54]  = 8'h3;
        test_receive_vector[55]  = 8'h3;
        test_receive_vector[56]  = 8'h3;
        test_receive_vector[57]  = 8'h4;
        test_receive_vector[58]  = 8'h3;
        test_receive_vector[59]  = 8'h5;
        test_receive_vector[60]  = 8'h3;
        test_receive_vector[61]  = 8'h6;
        test_receive_vector[62]  = 8'h3;
        test_receive_vector[63]  = 8'h7;
        test_receive_vector[64]  = 8'h4;
        test_receive_vector[65]  = 8'h0;
        test_receive_vector[66]  = 8'h4;
        test_receive_vector[67]  = 8'h1;
        test_receive_vector[68]  = 8'h4;
        test_receive_vector[69]  = 8'h2;
        test_receive_vector[70]  = 8'h4;
        test_receive_vector[71]  = 8'h3;
        test_receive_vector[72]  = 8'h4;
        test_receive_vector[73]  = 8'h4;
        test_receive_vector[74]  = 8'h4;
        test_receive_vector[75]  = 8'h5;
        test_receive_vector[76]  = 8'h4;
        test_receive_vector[77]  = 8'h6;
        test_receive_vector[78]  = 8'h4;
        test_receive_vector[79]  = 8'h7;
        test_receive_vector[80]  = 8'h5;
        test_receive_vector[81]  = 8'h0;
        test_receive_vector[82]  = 8'h5;
        test_receive_vector[83]  = 8'h1;
        test_receive_vector[84]  = 8'h5;
        test_receive_vector[85]  = 8'h2;
        test_receive_vector[86]  = 8'h5;
        test_receive_vector[87]  = 8'h3;
        test_receive_vector[88]  = 8'h5;
        test_receive_vector[89]  = 8'h4;
        test_receive_vector[90]  = 8'h5;
        test_receive_vector[91]  = 8'h5;
        test_receive_vector[92]  = 8'h5;
        test_receive_vector[93]  = 8'h6;
        test_receive_vector[94]  = 8'h5;
        test_receive_vector[95]  = 8'h7;
        test_receive_vector[96]  = 8'h6;
        test_receive_vector[97]  = 8'h0;
        test_receive_vector[98]  = 8'h6;
        test_receive_vector[99]  = 8'h1;
        test_receive_vector[100]  = 8'h6;
        test_receive_vector[101]  = 8'h2;
        test_receive_vector[102]  = 8'h6;
        test_receive_vector[103]  = 8'h3;
        test_receive_vector[104]  = 8'h6;
        test_receive_vector[105]  = 8'h4;
        test_receive_vector[106]  = 8'h6;
        test_receive_vector[107]  = 8'h5;
        test_receive_vector[108]  = 8'h6;
        test_receive_vector[109]  = 8'h6;
        test_receive_vector[110]  = 8'h6;
        test_receive_vector[111]  = 8'h7;
        test_receive_vector[112]  = 8'h7;
        test_receive_vector[113]  = 8'h0;
        test_receive_vector[114]  = 8'h7;
        test_receive_vector[115]  = 8'h1;
        test_receive_vector[116]  = 8'h7;
        test_receive_vector[117]  = 8'h2;
        test_receive_vector[118]  = 8'h7;
        test_receive_vector[119]  = 8'h3;
        test_receive_vector[120]  = 8'h7;
        test_receive_vector[121]  = 8'h4;
        test_receive_vector[122]  = 8'h7;
        test_receive_vector[123]  = 8'h5;
        test_receive_vector[124]  = 8'h7;
        test_receive_vector[125]  = 8'h6;
        test_receive_vector[126]  = 8'h7;
        test_receive_vector[127]  = 8'h7;
        test_receive_vector[128]  = 8'h8;
        test_receive_vector[129]  = 8'h0;
        test_receive_vector[130]  = 8'h8;
        test_receive_vector[131]  = 8'h1;
        test_receive_vector[132]  = 8'h8;
        test_receive_vector[133]  = 8'h2;
        test_receive_vector[134]  = 8'h8;
        test_receive_vector[135]  = 8'h3;
        test_receive_vector[136]  = 8'h8;
        test_receive_vector[137]  = 8'h4;
        test_receive_vector[138]  = 8'h8;
        test_receive_vector[139]  = 8'h5;
        test_receive_vector[140]  = 8'h8;
        test_receive_vector[141]  = 8'h6;
        test_receive_vector[142]  = 8'h8;
        test_receive_vector[143]  = 8'h7;
        test_receive_vector[144]  = 8'h9;
        test_receive_vector[145]  = 8'h0;
        test_receive_vector[146]  = 8'h9;
        test_receive_vector[147]  = 8'h1;
        test_receive_vector[148]  = 8'h9;
        test_receive_vector[149]  = 8'h2;
        test_receive_vector[150]  = 8'h9;
        test_receive_vector[151]  = 8'h3;
        test_receive_vector[152]  = 8'h9;
        test_receive_vector[153]  = 8'h4;
        test_receive_vector[154]  = 8'h9;
        test_receive_vector[155]  = 8'h5;
        test_receive_vector[156]  = 8'h9;
        test_receive_vector[157]  = 8'h6;
        test_receive_vector[158]  = 8'h9;
        test_receive_vector[159]  = 8'h7;
        test_receive_vector[160]  = 8'ha;
        test_receive_vector[161]  = 8'h0;
        test_receive_vector[162]  = 8'ha;
        test_receive_vector[163]  = 8'h1;
        test_receive_vector[164]  = 8'ha;
        test_receive_vector[165]  = 8'h2;
        test_receive_vector[166]  = 8'ha;
        test_receive_vector[167]  = 8'h3;
        test_receive_vector[168]  = 8'ha;
        test_receive_vector[169]  = 8'h4;
        test_receive_vector[170]  = 8'ha;
        test_receive_vector[171]  = 8'h5;
        test_receive_vector[172]  = 8'ha;
        test_receive_vector[173]  = 8'h6;
        test_receive_vector[174]  = 8'ha;
        test_receive_vector[175]  = 8'h7;
        test_receive_vector[176]  = 8'hb;
        test_receive_vector[177]  = 8'h0;
        test_receive_vector[178]  = 8'hb;
        test_receive_vector[179]  = 8'h1;
        test_receive_vector[180]  = 8'hb;
        test_receive_vector[181]  = 8'h2;
        test_receive_vector[182]  = 8'hb;
        test_receive_vector[183]  = 8'h3;
        test_receive_vector[184]  = 8'hb;
        test_receive_vector[185]  = 8'h4;
        test_receive_vector[186]  = 8'hb;
        test_receive_vector[187]  = 8'h5;
        test_receive_vector[188]  = 8'hb;
        test_receive_vector[189]  = 8'h6;
        test_receive_vector[190]  = 8'hb;
        test_receive_vector[191]  = 8'h7;
        test_receive_vector[192]  = 8'hc;
        test_receive_vector[193]  = 8'h0;
        test_receive_vector[194]  = 8'hc;
        test_receive_vector[195]  = 8'h1;
        test_receive_vector[196]  = 8'hc;
        test_receive_vector[197]  = 8'h2;
        test_receive_vector[198]  = 8'hc;
        test_receive_vector[199]  = 8'h3;
        test_receive_vector[200]  = 8'hc;
        test_receive_vector[201]  = 8'h4;
        test_receive_vector[202]  = 8'hc;
        test_receive_vector[203]  = 8'h5;
        test_receive_vector[204]  = 8'hc;
        test_receive_vector[205]  = 8'h6;
        test_receive_vector[206]  = 8'hc;
        test_receive_vector[207]  = 8'h7;
        test_receive_vector[208]  = 8'hd;
        test_receive_vector[209]  = 8'h0;
        test_receive_vector[210]  = 8'hd;
        test_receive_vector[211]  = 8'h1;
        test_receive_vector[212]  = 8'hd;
        test_receive_vector[213]  = 8'h2;
        test_receive_vector[214]  = 8'hd;
        test_receive_vector[215]  = 8'h3;
        test_receive_vector[216]  = 8'hd;
        test_receive_vector[217]  = 8'h4;
        test_receive_vector[218]  = 8'hd;
        test_receive_vector[219]  = 8'h5;
        test_receive_vector[220]  = 8'hd;
        test_receive_vector[221]  = 8'h6;
        test_receive_vector[222]  = 8'hd;
        test_receive_vector[223]  = 8'h7;
        test_receive_vector[224]  = 8'he;
        test_receive_vector[225]  = 8'h0;
        test_receive_vector[226]  = 8'he;
        test_receive_vector[227]  = 8'h1;
        test_receive_vector[228]  = 8'he;
        test_receive_vector[229]  = 8'h2;
        test_receive_vector[230]  = 8'he;
        test_receive_vector[231]  = 8'h3;
        test_receive_vector[232]  = 8'he;
        test_receive_vector[233]  = 8'h4;
        test_receive_vector[234]  = 8'he;
        test_receive_vector[235]  = 8'h5;
        test_receive_vector[236]  = 8'he;
        test_receive_vector[237]  = 8'h6;
        test_receive_vector[238]  = 8'he;
        test_receive_vector[239]  = 8'h7;
        test_receive_vector[240]  = 8'hf;
        test_receive_vector[241]  = 8'h0;
        test_receive_vector[242]  = 8'hf;
        test_receive_vector[243]  = 8'h1;
        test_receive_vector[244]  = 8'hf;
        test_receive_vector[245]  = 8'h2;
        test_receive_vector[246]  = 8'hf;
        test_receive_vector[247]  = 8'h3;
        test_receive_vector[248]  = 8'hf;
        test_receive_vector[249]  = 8'h4;
        test_receive_vector[250]  = 8'hf;
        test_receive_vector[251]  = 8'h5;
        test_receive_vector[252]  = 8'hf;
        test_receive_vector[253]  = 8'h6;
        test_receive_vector[254]  = 8'hf;
        test_receive_vector[255]  = 8'h7;
        test_receive_vector[256]  = 8'h10;
        test_receive_vector[257]  = 8'h0;
        test_receive_vector[258]  = 8'h10;
        test_receive_vector[259]  = 8'h1;
        test_receive_vector[260]  = 8'h10;
        test_receive_vector[261]  = 8'h2;
        test_receive_vector[262]  = 8'h10;
        test_receive_vector[263]  = 8'h3;
        test_receive_vector[264]  = 8'h10;
        test_receive_vector[265]  = 8'h4;
        test_receive_vector[266]  = 8'h10;
        test_receive_vector[267]  = 8'h5;
        test_receive_vector[268]  = 8'h10;
        test_receive_vector[269]  = 8'h6;
        test_receive_vector[270]  = 8'h10;
        test_receive_vector[271]  = 8'h7;
        test_receive_vector[272]  = 8'h11;
        test_receive_vector[273]  = 8'h0;
        test_receive_vector[274]  = 8'h11;
        test_receive_vector[275]  = 8'h1;
        test_receive_vector[276]  = 8'h11;
        test_receive_vector[277]  = 8'h2;
        test_receive_vector[278]  = 8'h11;
        test_receive_vector[279]  = 8'h3;
        test_receive_vector[280]  = 8'h11;
        test_receive_vector[281]  = 8'h4;
        test_receive_vector[282]  = 8'h11;
        test_receive_vector[283]  = 8'h5;
        test_receive_vector[284]  = 8'h11;
        test_receive_vector[285]  = 8'h6;
        test_receive_vector[286]  = 8'h11;
        test_receive_vector[287]  = 8'h7;
        test_receive_vector[288]  = 8'h12;
        test_receive_vector[289]  = 8'h0;
        test_receive_vector[290]  = 8'h12;
        test_receive_vector[291]  = 8'h1;
        test_receive_vector[292]  = 8'h12;
        test_receive_vector[293]  = 8'h2;
        test_receive_vector[294]  = 8'h12;
        test_receive_vector[295]  = 8'h3;
        test_receive_vector[296]  = 8'h12;
        test_receive_vector[297]  = 8'h4;
        test_receive_vector[298]  = 8'h12;
        test_receive_vector[299]  = 8'h5;
        test_receive_vector[300]  = 8'h12;
        test_receive_vector[301]  = 8'h6;
        test_receive_vector[302]  = 8'h12;
        test_receive_vector[303]  = 8'h7;
        test_receive_vector[304]  = 8'h13;
        test_receive_vector[305]  = 8'h0;
        test_receive_vector[306]  = 8'h13;
        test_receive_vector[307]  = 8'h1;
        test_receive_vector[308]  = 8'h13;
        test_receive_vector[309]  = 8'h2;
        test_receive_vector[310]  = 8'h13;
        test_receive_vector[311]  = 8'h3;
        test_receive_vector[312]  = 8'h13;
        test_receive_vector[313]  = 8'h4;
        test_receive_vector[314]  = 8'h13;
        test_receive_vector[315]  = 8'h5;
        test_receive_vector[316]  = 8'h13;
        test_receive_vector[317]  = 8'h6;
        test_receive_vector[318]  = 8'h13;
        test_receive_vector[319]  = 8'h7;
        test_receive_vector[320]  = 8'h14;
        test_receive_vector[321]  = 8'h0;
        test_receive_vector[322]  = 8'h14;
        test_receive_vector[323]  = 8'h1;
        test_receive_vector[324]  = 8'h14;
        test_receive_vector[325]  = 8'h2;
        test_receive_vector[326]  = 8'h14;
        test_receive_vector[327]  = 8'h3;
        test_receive_vector[328]  = 8'h14;
        test_receive_vector[329]  = 8'h4;
        test_receive_vector[330]  = 8'h14;
        test_receive_vector[331]  = 8'h5;
        test_receive_vector[332]  = 8'h14;
        test_receive_vector[333]  = 8'h6;
        test_receive_vector[334]  = 8'h14;
        test_receive_vector[335]  = 8'h7;
        test_receive_vector[336]  = 8'h15;
        test_receive_vector[337]  = 8'h0;
        test_receive_vector[338]  = 8'h15;
        test_receive_vector[339]  = 8'h1;
        test_receive_vector[340]  = 8'h15;
        test_receive_vector[341]  = 8'h2;
        test_receive_vector[342]  = 8'h15;
        test_receive_vector[343]  = 8'h3;
        test_receive_vector[344]  = 8'h15;
        test_receive_vector[345]  = 8'h4;
        test_receive_vector[346]  = 8'h15;
        test_receive_vector[347]  = 8'h5;
        test_receive_vector[348]  = 8'h15;
        test_receive_vector[349]  = 8'h6;
        test_receive_vector[350]  = 8'h15;
        test_receive_vector[351]  = 8'h7;
        test_receive_vector[352]  = 8'h16;
        test_receive_vector[353]  = 8'h0;
        test_receive_vector[354]  = 8'h16;
        test_receive_vector[355]  = 8'h1;
        test_receive_vector[356]  = 8'h16;
        test_receive_vector[357]  = 8'h2;
        test_receive_vector[358]  = 8'h16;
        test_receive_vector[359]  = 8'h3;
        test_receive_vector[360]  = 8'h16;
        test_receive_vector[361]  = 8'h4;
        test_receive_vector[362]  = 8'h16;
        test_receive_vector[363]  = 8'h5;
        test_receive_vector[364]  = 8'h16;
        test_receive_vector[365]  = 8'h6;
        test_receive_vector[366]  = 8'h16;
        test_receive_vector[367]  = 8'h7;
        test_receive_vector[368]  = 8'h17;
        test_receive_vector[369]  = 8'h0;
        test_receive_vector[370]  = 8'h17;
        test_receive_vector[371]  = 8'h1;
        test_receive_vector[372]  = 8'h17;
        test_receive_vector[373]  = 8'h2;
        test_receive_vector[374]  = 8'h17;
        test_receive_vector[375]  = 8'h3;
        test_receive_vector[376]  = 8'h17;
        test_receive_vector[377]  = 8'h4;
        test_receive_vector[378]  = 8'h17;
        test_receive_vector[379]  = 8'h5;
        test_receive_vector[380]  = 8'h17;
        test_receive_vector[381]  = 8'h6;
        test_receive_vector[382]  = 8'h17;
        test_receive_vector[383]  = 8'h7;
    end
    // Outputs
    wire tx;
    wire [23:0] leds;

    // Instantiate the Unit Under Test (UUT)
    lights uut (
        .clk(clk),
        .rx(rx),
        .tx(tx),
        .leds(leds)
    );

    always #20 clk = ~clk;

    // Transmission loop
    initial begin
        // Wait 100 ns for global reset to finish and a little longer for good measure.
        #100;
        #1234;

        for (i=0; i<test_send_vector_len; i=i+1) begin
            $display("Send i: %d val: %x", i, test_send_vector[i]);
            xmit_byte(test_send_vector[i]);
            if ((i+1) % 3 == 0) @ (test_step_complete) test_step_complete = 0; // Wait for module to echo result back to us
            // Wait random time
            random_delay = $random % 1000000; // Up to 1 ms
            #(random_delay);
        end

        #1000000
        if (write_complete_received == 0)   $display("Test failed");
        else                                $display("Test passed");
        $stop;
    end
    
    // Receiver loop
    always begin
        for (j=0; j<test_receive_vector_len; j=j+1) begin
            recv_byte(received_byte);
            $display("Recv j: %d expect: %x val: %x", j, test_receive_vector[j], received_byte);
            if (received_byte != test_receive_vector[j]) $stop;
            if ((j+1) % 2 == 0) test_step_complete = 1;
        end

        write_complete_received = 1;
    end

    task xmit_byte();
        input [7:0] b;
        integer i;
        begin
            #8681 rx = 0; xmit = 1; // start bit

            for (i=0;i<8;i = i+1) begin
                #8681 rx = b[0]; xmit = 0; // 0
                b = {1'b0, b[7:1]};
            end

            #8681 rx = 1; // stop bit
        end
    endtask
    
    task recv_byte();
        output [7:0] b;
        integer i;
        begin
            b = 0;
            @ (negedge tx); // Wait for start bit
            recv = 1;
            #4340;          // Wait half a bit period to align sampling to middle of transition.
            // 8 times, wait a bit period and then sample the value, shifting in from left to right.
            for (i=0;i<8;i = i+1) begin
                b = {1'b0, b[7:1]};
                #8681 b[7] = tx; recv = 0;
            end
            #4340;          // Wait another half a bit period to give the stop bit some time to occur.
        end
    endtask
    
endmodule

